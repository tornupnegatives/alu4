

***********************************************************
* CDL produced by pvsBuildNetlist on Apr  4 18:27:50 2024 *
***********************************************************


*pvsViewList = auLvs schematic
*pvsStopList = ("auLvs")
*pvsSimName  = auLvs



*.EXPAND_ON_M_FACTOR
*.MEGA

*.GLOBAL
+  vdd!
+  gnd!




* IGNORE_DUP_WARN
.subckt gnd gnd!
*PVSCELL netlisted from basic gnd schematic
*.generic no
.ends gnd


* IGNORE_DUP_WARN
.subckt vdd vdd!
*PVSCELL netlisted from basic vdd schematic
*.generic no
.ends vdd


.subckt inv1 a y
*PVSCELL netlisted from std_cells inv1 schematic
  MNM1 y a gnd! gnd! nfet_01v8 m=1 l=150n w=520n
  MPM0 y a vdd! vdd! pfet_01v8 m=1 l=150n w=1.66u
.ends inv1


.subckt nor2 a b y
*PVSCELL netlisted from std_cells nor2 schematic
  MNM0 y a gnd! gnd! nfet_01v8 m=1 l=150n w=520n
  MNM1 y b gnd! gnd! nfet_01v8 m=1 l=150n w=520n
  MPM0 net1 a vdd! vdd! pfet_01v8 m=1 l=150n w=1.04u
  MPM1 y b net1 vdd! pfet_01v8 m=1 l=150n w=1.04u
.ends nor2


.subckt or2 a b y
*PVSCELL netlisted from std_cells or2 schematic
  XI1 inv1 $PINS a=net1 y=y
  XI0 nor2 $PINS a=a b=b y=net1
.ends or2


***********************************************************
*             Completed at Apr  4 18:27:50 2024           *
***********************************************************
