* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : and2                                         *
* Netlisted  : Thu Apr  4 22:31:21 2024                     *
* Pegasus Version: 21.32-s016 Wed Nov 9 21:23:04 PST 2022   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 R(res_generic_m1) met1_res met1(P) met1(N)
*.DEVTMPLT 1 R(res_generic_m2) met2_res met2(P) met2(N)
*.DEVTMPLT 2 R(res_generic_m3) met3_res met3(P) met3(N)
*.DEVTMPLT 3 R(res_generic_m4) met4_res met4(P) met4(N)
*.DEVTMPLT 4 R(res_generic_m5) met5_res met5(P) met5(N)
*.DEVTMPLT 5 R(RES_GENERIC_ND) diff_res np_term(P) np_term(N)
*.DEVTMPLT 6 R(RES_GENERIC_PD) diff_res pp_term(P) pp_term(N)
*.DEVTMPLT 7 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 8 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_6                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_6 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_7                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_7 1 2 3 4
** N=6 EP=4 FDC=1
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=7.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_8                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_8 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=7.8e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_9                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_9 1 2 3
** N=7 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=7.8e-07 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nand2                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nand2 vdd! gnd! a b y
** N=11 EP=5 FDC=4
X5 vdd! y a pfet_01v8_CDNS_6 $T=645 4680 1 180 $X=50 $Y=4500
X6 6 y b gnd! nfet_01v8_CDNS_7 $T=925 520 0 0 $X=810 $Y=370
X7 gnd! 6 a nfet_01v8_CDNS_8 $T=495 520 0 0 $X=90 $Y=370
X8 vdd! y b pfet_01v8_CDNS_9 $T=925 4680 0 0 $X=520 $Y=4500
.ends nand2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_12                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_12 1 2 3
** N=5 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=5.2e-07 $X=0 $Y=0 $dt=7
.ends nfet_01v8_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_13                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_13 1 2 3
** N=11 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1.66e-06 $X=0 $Y=0 $dt=8
.ends pfet_01v8_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv1 vdd! gnd! a y
** N=6 EP=4 FDC=2
X2 gnd! y a nfet_01v8_CDNS_12 $T=495 520 0 0 $X=90 $Y=370
X3 vdd! y a pfet_01v8_CDNS_13 $T=495 3800 0 0 $X=50 $Y=3620
.ends inv1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: and2                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt and2 ain bin gnd! vdd! yout
** N=6 EP=5 FDC=6
X2 vdd! gnd! ain bin 1 nand2 $T=0 0 0 0 $X=0 $Y=-260
X3 vdd! gnd! 1 yout inv1 $T=1475 0 0 0 $X=1475 $Y=-260
.ends and2
