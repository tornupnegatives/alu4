`timescale 1ns / 1ps

module not1(
    input a,
    output logic r
    );
    not i0(r,a);
endmodule
